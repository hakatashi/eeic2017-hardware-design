module mul4(result, A, B);
	output [7:0] result;
	input [3:0] A, B;
	assign result = A * B;
endmodule
