module sub4(result, A, B);
	output [4:0] result;
	input [3:0] A, B;
	assign result = A - B;
endmodule
